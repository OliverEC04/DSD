library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity my_gates is
	port
	( 
		-- inputs
		

		-- outputs
		
	);
end my_gates;

architecture my_gates_impl of my_gates is

	function my_xor

begin

end my_gates_impl;
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.ALL;
ENTITY hex_mux IS
	PORT (
		-- Input ports
		

		-- Output ports
		
	);
END hex_mux;

ARCHITECTURE hex_mux_impl OF hex_mux IS
BEGIN
	
END hex_mux_impl;
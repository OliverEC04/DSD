library verilog;
use verilog.vl_types.all;
entity four_bit_adder_tester_vlg_vec_tst is
end four_bit_adder_tester_vlg_vec_tst;
